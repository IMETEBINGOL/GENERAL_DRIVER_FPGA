localparam  CAC_SETTINGS_MEMORY_WIDTH           = 16;
localparam  CAC_SETTINGS_ROM_MEMORY_LENGTH      = 16;
localparam  CAC_SETTINGS_RAM_MEMORY_LENGTH      = 16;
localparam  CAC_UART_BAUDRATE                   = 115200;
localparam  CAC_UART_BITLEN                     = 8;
localparam  CAC_UART_BUFFER_WIDTH               = 8;
localparam  CAC_UART_BUFFER_DEPTH               = 16;
localparam  CAC_UART_ERRORNUM                   = 3;
localparam  CAC_BUFFER_WIDTH                    = 8;
localparam  CAC_SPI_PACKAGE_WIDTH               = 8;