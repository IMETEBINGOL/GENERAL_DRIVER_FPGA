`define SPI_WRITE   0'h01
`define SPI_READ    0'h02