localparam  COMMAND_INITIAL_STATE   = 0;
// UART RESET STATES
// ---
localparam  UART_RESET_PROCESS_0    = 1;
localparam  UART_RESET_PROCESS_1    = 2;
localparam  UART_RESET_PROCESS_2    = 3;
localparam  UART_RESET_PROCESS_3    = 4;
localparam  UART_RESET_PROCESS_4    = 5;
// ---
// SETTINGS WRITE STATES
// ---
localparam  UART_WRITEREG_PROCESS_0 = 1; 
localparam  UART_WRITEREG_PROCESS_1 = 2;
localparam  UART_WRITEREG_PROCESS_2 = 3;
localparam  UART_WRITEREG_PROCESS_3 = 4;
localparam  UART_WRITEREG_PROCESS_4 = 5;
localparam  UART_WRITEREG_PROCESS_5 = 6;
localparam  UART_WRITEREG_PROCESS_6 = 7;
localparam  UART_WRITEREG_PROCESS_7 = 8;
// ---
// SETTINGS READ STATES
// ---
localparam  UART_READREG_PROCESS_0  = 1;
localparam  UART_READREG_PROCESS_1  = 2;
localparam  UART_READREG_PROCESS_2  = 3;
localparam  UART_READREG_PROCESS_3  = 4;
localparam  UART_READREG_PROCESS_4  = 5;
// ---





