case (cmd_spi)
    `include "../COMMANDS/SPI_WRITE/spi_write.vh"
    `include "../COMMANDS/SPI_READ/spi_read.vh"
    `include "../COMMANDS/DEFAULT/default.vh"
endcase