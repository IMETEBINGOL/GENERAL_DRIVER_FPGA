`SPI_READ:
begin
    case (cmd_state)
        COMMAND_STATE_INITIAL:
        begin
            
        end
        COMMAND_READ_PROCESS_0:
        begin
            
        end
        COMMAND_READ_PROCESS_1:
        begin
            
        end
        COMMAND_READ_PROCESS_2:
        begin
            
        end 
        default:
        begin
            
        end 
    endcase
end