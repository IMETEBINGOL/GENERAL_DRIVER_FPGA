`define SPI_WRITE   8'h01
`define SPI_READ    8'h02