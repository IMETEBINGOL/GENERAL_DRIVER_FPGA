localparam  CAC_CLK_FREQUENCY   = 10_000_000;