`define UARTRST_OPCODE  8'h10
`define WRITEREG_OPCODE 8'h01
`define READREG_OPCODE  8'h02