localparam  MASTER_CLOCK_FREQUENCY   = 100_000_000;   