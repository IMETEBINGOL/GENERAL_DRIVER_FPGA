default:
begin
    state_reset();
end