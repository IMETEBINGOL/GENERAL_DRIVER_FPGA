case (command)
    `include "../COMMANDS/UARTRST/uartrst.vh"
    `include "../COMMANDS/WRITEREG/writereg.vh"
    `include "../COMMANDS/READREG/readreg.vh"
    `include "../COMMANDS/DEFAULT/default.vh"
endcase