default:
begin
    state   <= CMDREAD; 
end