assign rom_memory[0]        = rom_data_0;
assign rom_memory[1]        = rom_data_1;
assign rom_memory[2]        = rom_data_2;
assign rom_memory[3]        = rom_data_3;
assign rom_memory[4]        = rom_data_4;
assign rom_memory[5]        = rom_data_5;
assign rom_memory[6]        = rom_data_6;
assign rom_memory[7]        = rom_data_7;
assign rom_memory[8]        = rom_data_8;
assign rom_memory[9]        = rom_data_9;
assign rom_memory[10]       = rom_data_10;
assign rom_memory[11]       = rom_data_11;
assign rom_memory[12]       = rom_data_12;
assign rom_memory[13]       = rom_data_13;
assign rom_memory[14]       = rom_data_14;
assign rom_memory[15]       = rom_data_15;