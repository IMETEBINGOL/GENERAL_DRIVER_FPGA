ram_memory[0]   <= 32'b00000000000000000000000000000000;
ram_memory[1]   <= 32'b00000000000000000000000000000000;
ram_memory[2]   <= 32'b00000000000000000000000000000000;
ram_memory[3]   <= 32'b00000000000000000000000000000000;
ram_memory[4]   <= 32'b00000000000000000000000000000000;
ram_memory[5]   <= 32'b00000000000000000000000000000000;
ram_memory[6]   <= 32'b00000000000000000000000000000000;
ram_memory[7]   <= 32'b00000000000000000000000000000000;
ram_memory[8]   <= 32'b00000000000000000000000000000000;
ram_memory[9]   <= 32'b00000000000000000000000000000000;
ram_memory[10]  <= 32'b00000000000000000000000000000000;
ram_memory[11]  <= 32'b00000000000000000000000000000000;
ram_memory[12]  <= 32'b00000000000000000000000000000000;
ram_memory[13]  <= 32'b00000000000000000000000000000000;
ram_memory[14]  <= 32'b00000000000000000000000000000000;
ram_memory[15]  <= 32'b00000000000000000000000000000000;