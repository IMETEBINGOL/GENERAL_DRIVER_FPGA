localparam      COMMAND_STATE_INITIAL   = 0;
// SPI READ PARAMETER 
localparam      COMMAND_READ_PROCESS_0  = 1;
localparam      COMMAND_READ_PROCESS_1  = 2;
localparam      COMMAND_READ_PROCESS_2  = 3;
// SPI WRITE PARAMETER 
localparam      COMMAND_WRITE_PROCESS_0  = 1;
localparam      COMMAND_WRITE_PROCESS_1  = 2;
localparam      COMMAND_WRITE_PROCESS_2  = 3;
